library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity elevador is
  port (
    M, F1, F2, F3 : in  std_logic;
    ABRIR, TRAVA : out std_logic );
end entity;

architecture  rtl OF elevador IS

begin


end architecture;
