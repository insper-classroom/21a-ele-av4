library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mapaKarnaught is
  port (
    A,B,C,D  : in  std_logic;
    S0,S1,S2,S3 : out std_logic );
end entity;

architecture  rtl OF mapaKarnaught IS

begin


end architecture;
